`define no_of_transaction 100
`define DSIZE 8
`define ASIZE 4
