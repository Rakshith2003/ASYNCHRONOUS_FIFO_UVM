package asy_fifo_pkg;
  `include "uvm_pkg.sv"
  `include "uvm_macros.svh"
  `include "asy_fifo_write_seq_item.sv"
  `include "asy_fifo_read_seq_item.sv"
  `include "asy_fifo_write_sequence.sv"
  `include "asy_fifo_read_sequence.sv"
  `include "asy_fifo_write_sequencer.sv"
  `include "asy_fifo_read_sequencer.sv"
  `include "virtual_sequencer.sv"
  `include "virtual_sequence.sv"

  `include "asy_fifo_write_driver.sv"
  `include "asy_fifo_read_driver.sv"
  `include "asy_fifo_write_monitor.sv"
  `include "asy_fifo_read_monitor.sv"
  `include "asy_fifo_write_agent.sv"
  `include "asy_fifo_read_agent.sv"
  `include "asy_fifo_scoreboard.sv"
  `include "asy_fifo_subscriber.sv"
  `include "asy_fifo_environment.sv"

  `include "asy_fifo_test.sv"

  //`include"alu_coverage.sv"

endpackage
